----------------------------------------------------------------------------------
-- Company: Trinity College Dublin
-- Engineer: Faith Olopade
-- 
-- Create Date: 17.10.2022 22:35:00
-- Design Name: 
-- Module Name: CPU_ControlMemory_21364066 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity CPU_ControlMemory_21364066 is
    port (
        Address : in std_logic_vector (16 downto 0);
        NA : out std_logic_vector (16 downto 0); -- 34-50
        MS : out std_logic_vector (2 downto 0); -- 31-33
        MC : out std_logic; -- 30
        IL : out std_logic; -- 29
        PI : out std_logic; -- 28
        PL : out std_logic; -- 27
        TD : out std_logic_vector (3 downto 0); -- 23-26
        TA : out std_logic_vector (3 downto 0); -- 19-22
        TB : out std_logic_vector (3 downto 0); -- 15-18
        MB : out std_logic; -- 14
        FS : out std_logic_vector (4 downto 0); -- 09-13
        MD : out std_logic; -- 08
        RW : out std_logic; -- 07
        MM : out std_logic; -- 06
        MW : out std_logic; -- 05
        RV : out std_logic; -- 04
        RC : out std_logic; -- 03
        RN : out std_logic; -- 02
        RZ : out std_logic; -- 01
        FL : out std_logic -- 00
        );
end CPU_ControlMemory_21364066;

architecture Behavioral of CPU_ControlMemory_21364066 is

    -- we use the least significant 7 bit of the Address - array(0 to 127)
type ROM_array is array(0 to 127) of std_logic_vector (50 downto 0);
signal ROM : ROM_array :=(
    --00 to 15--
--|50 34|33 31|30| 29| 28| 27|26 23|22 19|18 15| 14|13 09| 08| 07| 06| 05| 04| 03| 02| 01| 00| Control Mem
--| Next Address | MS |MC| IL| PI| PL| TD | TA | TB | MB| FS | MD| RW| MM| MW| RV| RC| RN| RZ| FL| Address      --INITIALIZE--
"00000000001000010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 0
"00000000001000011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 1
"00000000001000100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 2
"00000000001000101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 3
"00000000001000110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 4
"00000000001000111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 5
"00000000001001000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 6
"00000000001001001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 7
"00000000001001010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 8
"00000000001001011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 9
"00000000001001100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 10
"00000000001001101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 11
"00000000001001110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 12
"00000000001001111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 13
"00000000001010000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 14
"00000000001010001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 15

--16 to 31
--|50 34|33 31|30| 29| 28| 27|26 23|22 19|18 15| 14|13 09| 08| 07| 06| 05| 04| 03| 02| 01| 00| Control Mem
--| Next Address | MS |MC| IL| PI| PL| TD | TA | TB | MB| FS | MD| RW| MM| MW| RV| RC| RN| RZ| FL| Address
"00000000001010010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 16
"00000000001010011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 17
"00000000001010100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 18
"00000000001010101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 19
"00000000001010110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 20
"00000000001010111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 21
"00000000001011000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 22
"00000000001011001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 23
"00000000001011010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 24
"00000000001011011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 25
"00000000001011100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 26
"00000000001011101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 27
"00000000001011110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 28
"00000000001011111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 29
"00000000001100000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 30
"00000000001100001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 31

--32 to 47
--|50 34|33 31|30| 29| 28| 27|26 23|22 19|18 15| 14|13 09| 08| 07| 06| 05| 04| 03| 02| 01| 00| Control Mem
--| Next Address | MS |MC| IL| PI| PL| TD | TA | TB | MB| FS | MD| RW| MM| MW| RV| RC| RN| RZ| FL| Address
"00000000001100010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 32
"00000000001100011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 33
"00000000001100100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 34
"00000000001100101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 35
"00000000001100110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 36
"00000000001100111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 37
"00000000001101000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 38
"00000000001101001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 39 
"00000000001101010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 40
"00000000001101011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 41
"00000000001101100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 42
"00000000001101101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 43
"00000000001101110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 44
"00000000001101111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 45
"00000000001110000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 46
"00000000001110001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 47

--48 to 63
--|50 34|33 31|30| 29| 28| 27|26 23|22 19|18 15| 14|13 09| 08| 07| 06| 05| 04| 03| 02| 01| 00| Control Mem
--| Next Address | MS |MC| IL| PI| PL| TD | TA | TB | MB| FS | MD| RW| MM| MW| RV| RC| RN| RZ| FL| Address
"00000000001110010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 48
"00000000001110011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 49
"00000000001110100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 50
"00000000001110101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 51
"00000000001110110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 52
"00000000001110111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 53
"00000000001111000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 54
"00000000001111001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 55
"00000000001111010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 56
"00000000001111011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 57
"00000000001111100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 58
"00000000001111101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 59
"00000000001111110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 60
"00000000001111111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 61
"00000000010000000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 62
"00000000010000001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 63

--64 to 79
--|50 34|33 31|30| 29| 28| 27|26 23|22 19|18 15| 14|13 09| 08| 07| 06| 05| 04| 03| 02| 01| 00| Control Mem
--| Next Address | MS |MC| IL| PI| PL| TD | TA | TB | MB| FS | MD| RW| MM| MW| RV| RC| RN| RZ| FL| Address
"00000000010000010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 64
"00000000010000011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 65
"00000000010000100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 66
"00000000010000101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 67
"00000000010000110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 68
"00000000010000111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 69
"00000000010001000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 70
"00000000010001001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 71
"00000000010001010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 72
"00000000010001011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 73
"00000000010001100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 74
"00000000010001101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 75
"00000000010001110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 76
"00000000010001111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 77
"00000000010010000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 78
"00000000010010001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 79

--80 to 95
--|50 34|33 31|30| 29| 28| 27|26 23|22 19|18 15| 14|13 09| 08| 07| 06| 05| 04| 03| 02| 01| 00| Control Mem
--| Next Address | MS |MC| IL| PI| PL| TD | TA | TB | MB| FS | MD| RW| MM| MW| RV| RC| RN| RZ| FL| Address
"00000000010010010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 80
"00000000010010011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 81
"00000000010010100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 82
"00000000010010101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 83
"00000000010010110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 84
"00000000010010111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 85
"00000000010011000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 86
"00000000010011001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 87
"00000000010011010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 88
"00000000010011011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 89
"00000000010011100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 90
"00000000010011101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 91
"00000000010011110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 92
"00000000010011111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 93
"00000000010100000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 94
"00000000010100001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 95

--96 to 111
--|50 34|33 31|30| 29| 28| 27|26 23|22 19|18 15| 14|13 09| 08| 07| 06| 05| 04| 03| 02| 01| 00| Control Mem
--| Next Address | MS |MC| IL| PI| PL| TD | TA | TB | MB| FS | MD| RW| MM| MW| RV| RC| RN| RZ| FL| Address
"00000000010100010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 96
"00000000010100011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 97
"00000000010100100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 98
"00000000010100101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 99
"00000000010100110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 100
"00000000010100111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 101
"00000000010101000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 102
"00000000010101001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 103
"00000000010101010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 104
"00000000010101011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 105
"00000000010101100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 106
"00000000010101101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 107
"00000000010101110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 108
"00000000010101111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 109
"00000000010110000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 110
"00000000010110001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 111

--112 to 127--
--|50 34|33 31|30| 29| 28| 27|26 23|22 19|18 15| 14|13 09| 08| 07| 06| 05| 04| 03| 02| 01| 00| Control Mem
--| Next Address | MS |MC| IL| PI| PL| TD | TA | TB | MB| FS | MD| RW| MM| MW| RV| RC| RN| RZ| FL| Address
"00000000010110010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 112
"00000000010110011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 113
"00000000010110100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 114
"00000000010110101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 115
"00000000010110110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 116
"00000000010110111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 117
"00000000010111000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 118
"00000000010111001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 119
"00000000010111010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 120
"00000000010111011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 121
"00000000010111100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 122
"00000000010111101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 123
"00000000010111110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 124
"00000000010111111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 125
"00000000011000000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- Next Address = Last 2 ID + 126
"00000000011000001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'  -- Next Address = Last 2 ID + 127
);

signal content_at_address : std_logic_vector (50 downto 0);

begin
    content_at_address <= ROM(to_integer(unsigned(Address(6 downto 0)))) after 2ns;
    
    NA <= content_at_address(50 downto 34); -- 34-50
    MS <= content_at_address(33 downto 31); -- 31-33
    MC <= content_at_address(30); -- 30
    IL <= content_at_address(29); -- 29
    PI <= content_at_address(28); -- 28
    PL <= content_at_address(27); -- 27
    TD <= content_at_address(26 downto 23); -- 23-26
    TA <= content_at_address(22 downto 19); -- 19-22
    TB <= content_at_address(18 downto 15); -- 15-18
    MB <= content_at_address(14); -- 14
    FS <= content_at_address(13 downto 9); -- 09-13
    MD <= content_at_address(8); -- 08
    RW <= content_at_address(7); -- 07
    MM <= content_at_address(6); -- 06
    MW <= content_at_address(5); -- 05
    RV <= content_at_address(4); -- 04
    RC <= content_at_address(3); -- 03
    RN <= content_at_address(2); -- 02
    RZ <= content_at_address(1); -- 01
    FL <= content_at_address(0); -- 00
    
end Behavioral;
