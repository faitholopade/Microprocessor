------------------------------------------------------------------------------------
---- Company: Trinity College architecture
---- Engineer: Faith Olopade
---- 
---- Create Date: 17.10.2022 23:12:00
---- Design Name: 
---- Module Name: CPU_DFlipFlop_21364066_TB - Sim
---- Project Name: 
---- Target Devices: 
---- Tool Versions: 
---- Description: 
---- 
---- Dependencies: 
---- 
---- Revision:
---- Revision 0.01 - File Created
---- Additional Comments:
---- 
------------------------------------------------------------------------------------


--library IEEE;
--use IEEE.STD_LOGIC_1164.ALL;

---- Uncomment the following library declaration if using
---- arithmetic functions with Signed or Unsigned values
----use IEEE.NUMERIC_STD.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx leaf cells in this code.
----library UNISIM;
----use UNISIM.VComponents.all;

--entity CPU_DFlipFlop_21364066_TB is
----  Port ( ); We don't need ports
--end CPU_DFlipFlop_21364066_TB;

--architecture Sim of CPU_DFlipFlop_21364066_TB is
---- Component Declaration for the Unit Under Test (UUT)

--component CPU_DFlipFlop_21364066
--port ( 
--      );
--end component;

----Inputs
--    signal 
----Outputs
--    signal 

    
--begin
--	-- Instantiate the Unit Under Test (UUT)
	
--   uut: CPU_DFlipFlop_21364066 port map (
          
--        );

        
--   stim_proc: process

--   begin

--   end process;
--end Sim;