    In00_TB <= "00000001010001011111110101100010";
    In01_TB <= "00000001010001011111110101100011";
    In02_TB <= "00000001010001011111110101100100";
    In03_TB <= "00000001010001011111110101100101";
    In04_TB <= "00000001010001011111110101100110";
    In05_TB <= "00000001010001011111110101100111";
    In06_TB <= "00000001010001011111110101101000";
    In07_TB <= "00000001010001011111110101101001";
    In08_TB <= "00000001010001011111110101101010";
    In09_TB <= "00000001010001011111110101101011";
    In10_TB <= "00000001010001011111110101101100";
    In11_TB <= "00000001010001011111110101101101";
    In12_TB <= "00000001010001011111110101101110";
    In13_TB <= "00000001010001011111110101101111";
    In14_TB <= "00000001010001011111110101110000";
    In15_TB <= "00000001010001011111110101110001";
    In16_TB <= "00000001010001011111110101110010";
    In17_TB <= "00000001010001011111110101110011";
    In18_TB <= "00000001010001011111110101110100"; 
    In19_TB <= "00000001010001011111110101110101";
    In20_TB <= "00000001010001011111110101110110";
    In21_TB <= "00000001010001011111110101110111";
    In22_TB <= "00000001010001011111110101111000";
    In23_TB <= "00000001010001011111110101111001";
    In24_TB <= "00000001010001011111110101111010";
    In25_TB <= "00000001010001011111110101111011";
    In26_TB <= "00000001010001011111110101111100";
    In27_TB <= "00000001010001011111110101111101";
    In28_TB <= "00000001010001011111110101111110";
    In29_TB <= "00000001010001011111110101111111";
    In30_TB <= "00000001010001011111110110000000";
    In31_TB <= "00000001010001011111110110000001";